module rom_case(out, address);
	output reg [31:0] out;
	input  [15:0] address; // address- 16 deep memory  
	always @(address) begin
		case (address)
			16'h0000:  out = 32'b11010010100000000000000000100001; // MOVZ X1, 1
			16'h0004:  out = 32'b11010010100000000000000001000010; // MOVZ X2, 2
			16'h0008:  out = 32'b10001011000000100000000000100100; // ADD X4, X1, X2
			16'h000C:  out = 32'b11111000000000010000001111100100; // STUR X4, [XZR, 16]
			16'h000F:  out = 32'b11111000010000010000001111100101; // LDUR X5, [XZR, 16]
			16'h0010:  out = 32'b10010100000000000000000000001010; // BL 10
			16'h0014:  out = 32'b10110101000000000000000000100010; // CBNZ X2, 1
			16'h0018:  out = 32'b00010100000000000000000000000001; // B 1
			16'h001C:  out = 32'b00010111111111111111111111111001; // B -7
			16'h0020:  out = 32'b10110100000000000000000001100001; // CBZ X1, 3
			16'h0024:  out = 32'b11101011000000100000000000111111; // SUBS XZR, X1, X2
			16'h0028:  out = 32'b01010100000000000000000000100011; // B.LO 1
			16'h002C:  out = 32'b11111000000000001000001111100001; // STUR X1, [XZR, 8]
			16'h0030:  out = 32'b11111000010000001000001111100110; // LDUR X6, [XZR, 8]
			16'h0034:  out = 32'b11010010000000000000010011100111; // EORI X7, X7, 1
			16'h0038:  out = 32'b00010111111111111111111111111110; // B -2
			16'h003C:  out = 32'b10010001000000000000100000100001; // ADDI X1, X1, 2
			16'h0040:  out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
			16'h0044:  out = 32'b11010110000000000000001111000000; // BR X30
			default: out=32'hD60003E0; //BR XZR
		endcase
	end
endmodule
